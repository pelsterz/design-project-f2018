module NESController(

);


	
endmodule

	