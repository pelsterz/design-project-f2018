module SPIReader(
	input logic _c,
	input logic _l,
	input logic [7:0] d,
	output logic [3:0] move
);

